library verilog;
use verilog.vl_types.all;
entity corners_tb is
    generic(
        WIDTH           : integer := 320;
        HEIGTH          : integer := 240
    );
end corners_tb;
