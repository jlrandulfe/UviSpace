library verilog;
use verilog.vl_types.all;
entity erosion_tb is
end erosion_tb;
