library verilog;
use verilog.vl_types.all;
entity convolution_tb is
    generic(
        WIDTH           : integer := 8;
        HEIGHT          : integer := 8
    );
end convolution_tb;
