library verilog;
use verilog.vl_types.all;
entity sram_controller_tb is
end sram_controller_tb;
