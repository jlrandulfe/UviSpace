library verilog;
use verilog.vl_types.all;
entity connected_tb is
    generic(
        WIDTH           : integer := 160;
        HEIGHT          : integer := 120
    );
end connected_tb;
