library verilog;
use verilog.vl_types.all;
entity convolution3s_tb is
end convolution3s_tb;
